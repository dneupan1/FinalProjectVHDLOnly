-- unnamed.vhd

-- Generated using ACDS version 21.1 850

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unnamed is
	port (
		lcd_clk_clk        : out std_logic;        --      lcd_clk.clk
		ref_clk_clk        : in  std_logic := '0'; --      ref_clk.clk
		ref_reset_reset    : in  std_logic := '0'; --    ref_reset.reset
		reset_source_reset : out std_logic;        -- reset_source.reset
		vga_clk_clk        : out std_logic;        --      vga_clk.clk
		video_in_clk_clk   : out std_logic         -- video_in_clk.clk
	);
end entity unnamed;

architecture rtl of unnamed is
	component unnamed_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			video_in_clk_clk   : out std_logic;        -- clk
			vga_clk_clk        : out std_logic;        -- clk
			lcd_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component unnamed_video_pll_0;

begin

	video_pll_0 : component unnamed_video_pll_0
		port map (
			ref_clk_clk        => ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => ref_reset_reset,    --    ref_reset.reset
			video_in_clk_clk   => video_in_clk_clk,   -- video_in_clk.clk
			vga_clk_clk        => vga_clk_clk,        --      vga_clk.clk
			lcd_clk_clk        => lcd_clk_clk,        --      lcd_clk.clk
			reset_source_reset => reset_source_reset  -- reset_source.reset
		);

end architecture rtl; -- of unnamed
